LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 3, 18, 9, 7, 2, 14, 8, 8, 0, 0, 0, 10, 12, 2, 2, 
		7, 17, 8, 6, 7, 71, 0, 2, 0, 21, 0, 0, 7, 15, 8, 
		0, 33, 11, 10, 7, 32, 0, 0, 0, 49, 0, 0, 0, 0, 40, 
		0, 55, 0, 10, 4, 7, 11, 0, 0, 23, 0, 0, 0, 0, 42, 
		0, 45, 0, 0, 39, 0, 0, 0, 0, 29, 0, 0, 12, 0, 0, 
		0, 46, 0, 0, 111, 0, 20, 0, 0, 96, 0, 0, 8, 0, 0, 
		0, 27, 0, 0, 72, 38, 9, 0, 0, 96, 0, 0, 0, 13, 0, 
		0, 12, 0, 2, 0, 56, 0, 0, 0, 65, 0, 0, 9, 8, 0, 
		0, 5, 0, 49, 0, 0, 0, 16, 9, 0, 23, 0, 21, 38, 10, 
		14, 0, 0, 38, 0, 0, 6, 22, 0, 0, 0, 0, 39, 30, 0, 
		89, 0, 0, 88, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
		21, 30, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 7, 12, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 4, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 
		1, 2, 2, 0, 6, 0, 0, 0, 0, 8, 0, 0, 11, 20, 0, 
		0, 47, 0, 0, 2, 13, 0, 0, 7, 38, 0, 0, 0, 25, 19, 
		0, 65, 3, 6, 0, 21, 0, 0, 0, 81, 0, 0, 0, 0, 75, 
		0, 22, 0, 81, 0, 0, 0, 0, 0, 96, 0, 0, 0, 0, 29, 
		0, 0, 0, 0, 60, 0, 0, 0, 0, 150, 0, 0, 12, 0, 0, 
		0, 0, 13, 0, 61, 28, 0, 0, 0, 118, 0, 0, 0, 8, 0, 
		0, 0, 0, 0, 50, 54, 0, 0, 0, 66, 0, 0, 22, 0, 0, 
		0, 0, 0, 25, 0, 21, 0, 0, 34, 0, 17, 0, 17, 18, 0, 
		0, 0, 0, 53, 0, 0, 36, 0, 0, 0, 0, 4, 39, 32, 0, 
		49, 0, 0, 129, 0, 0, 20, 0, 0, 0, 1, 0, 0, 5, 0, 
		73, 30, 0, 69, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 64, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 123, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
		0, 0, 0, 3, 0, 7, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 11, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 4, 49, 13, 0, 0, 5, 9, 0, 
		21, 39, 0, 0, 0, 28, 42, 22, 0, 0, 0, 0, 0, 0, 3, 
		0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 4, 0, 19, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 6, 63, 8, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
		0, 0, 5, 18, 5, 0, 4, 0, 0, 0, 9, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 16, 23, 7, 0, 19, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 38, 8, 0, 0, 1, 14, 43, 5, 0, 0, 
		12, 0, 3, 0, 0, 0, 0, 0, 0, 32, 51, 15, 0, 0, 0, 
		23, 0, 13, 0, 0, 0, 0, 34, 17, 11, 0, 0, 0, 17, 29, 
		20, 31, 0, 0, 75, 81, 40, 36, 19, 6, 0, 0, 0, 0, 0, 
		0, 3, 0, 5, 68, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
		0, 0, 0, 98, 23, 0, 0, 0, 0, 0, 0, 3, 5, 0, 17, 
		0, 0, 1, 47, 14, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		62, 63, 63, 63, 62, 62, 66, 69, 64, 61, 56, 57, 53, 50, 46, 
		58, 66, 66, 65, 65, 76, 56, 65, 56, 36, 22, 24, 41, 48, 49, 
		60, 72, 67, 65, 71, 109, 44, 27, 9, 54, 34, 20, 14, 24, 50, 
		4, 41, 64, 69, 65, 54, 41, 14, 20, 65, 41, 35, 11, 0, 48, 
		9, 62, 51, 67, 70, 60, 49, 18, 19, 39, 44, 13, 21, 0, 20, 
		35, 80, 47, 79, 117, 66, 58, 23, 5, 78, 65, 17, 31, 12, 0, 
		20, 83, 46, 47, 90, 77, 92, 47, 13, 106, 44, 14, 23, 25, 13, 
		44, 62, 21, 43, 57, 112, 72, 60, 18, 96, 49, 17, 28, 44, 25, 
		65, 84, 18, 55, 44, 65, 33, 37, 31, 65, 51, 21, 21, 27, 46, 
		90, 84, 24, 65, 24, 37, 49, 51, 36, 47, 25, 0, 21, 69, 65, 
		107, 85, 38, 91, 37, 18, 88, 86, 24, 13, 0, 0, 21, 45, 31, 
		87, 92, 44, 153, 108, 25, 36, 28, 3, 7, 8, 14, 9, 15, 9, 
		5, 67, 77, 145, 16, 7, 6, 6, 3, 2, 6, 10, 21, 19, 15, 
		0, 5, 89, 99, 10, 14, 3, 3, 6, 9, 15, 15, 7, 14, 34, 
		2, 3, 20, 38, 9, 14, 16, 8, 11, 12, 4, 4, 16, 23, 0, 
		
		98, 100, 101, 103, 98, 92, 109, 115, 100, 80, 70, 73, 82, 93, 90, 
		98, 103, 104, 106, 98, 54, 102, 81, 72, 17, 9, 18, 35, 63, 83, 
		66, 69, 100, 109, 104, 82, 71, 40, 14, 0, 29, 25, 26, 30, 60, 
		50, 0, 99, 94, 78, 43, 32, 31, 15, 6, 49, 32, 30, 26, 30, 
		46, 0, 105, 50, 28, 44, 57, 39, 23, 0, 32, 46, 13, 26, 18, 
		43, 14, 114, 69, 21, 67, 48, 44, 31, 0, 57, 54, 14, 21, 19, 
		46, 19, 75, 99, 12, 7, 44, 42, 50, 0, 59, 32, 6, 3, 39, 
		33, 25, 37, 56, 25, 7, 73, 38, 51, 2, 47, 40, 6, 33, 75, 
		26, 2, 45, 2, 37, 43, 47, 12, 14, 39, 29, 55, 15, 42, 72, 
		25, 14, 49, 0, 50, 28, 7, 17, 30, 49, 42, 8, 0, 44, 81, 
		0, 15, 51, 0, 26, 4, 0, 18, 33, 0, 0, 0, 0, 0, 0, 
		0, 0, 35, 0, 55, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 8, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 19, 0, 4, 0, 19, 17, 0, 0, 0, 
		16, 0, 0, 0, 0, 0, 32, 8, 0, 0, 49, 31, 53, 0, 0, 
		88, 0, 0, 0, 9, 0, 24, 31, 25, 0, 69, 25, 41, 33, 0, 
		81, 1, 40, 0, 18, 40, 72, 55, 42, 0, 35, 68, 15, 45, 0, 
		76, 24, 54, 21, 0, 30, 74, 48, 78, 0, 90, 69, 1, 33, 32, 
		66, 89, 6, 40, 0, 0, 47, 58, 75, 0, 92, 57, 13, 1, 45, 
		67, 69, 41, 25, 0, 0, 107, 36, 46, 0, 64, 66, 0, 23, 23, 
		84, 38, 116, 0, 39, 12, 35, 32, 0, 52, 0, 63, 0, 0, 1, 
		48, 43, 124, 0, 60, 16, 0, 53, 46, 19, 56, 1, 0, 0, 2, 
		0, 41, 117, 0, 128, 52, 0, 52, 77, 42, 3, 5, 14, 0, 14, 
		0, 2, 49, 0, 163, 74, 33, 34, 38, 26, 29, 31, 35, 41, 46, 
		68, 0, 0, 89, 120, 37, 44, 37, 36, 31, 30, 34, 44, 36, 30, 
		69, 41, 0, 121, 51, 32, 52, 40, 31, 35, 44, 42, 49, 22, 80, 
		83, 46, 46, 36, 44, 22, 30, 37, 32, 44, 57, 35, 8, 79, 92, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 9, 12, 0, 0, 
		9, 0, 0, 0, 0, 0, 0, 5, 7, 0, 8, 4, 15, 15, 0, 
		36, 0, 0, 0, 0, 0, 4, 13, 16, 0, 0, 14, 0, 10, 0, 
		68, 13, 0, 0, 0, 6, 0, 0, 13, 0, 27, 30, 1, 11, 13, 
		64, 30, 0, 0, 0, 0, 0, 10, 14, 0, 36, 25, 12, 3, 6, 
		61, 27, 29, 0, 0, 0, 33, 13, 6, 0, 14, 25, 6, 0, 0, 
		61, 41, 73, 0, 0, 6, 3, 0, 0, 0, 0, 24, 3, 0, 0, 
		29, 35, 57, 15, 31, 15, 0, 0, 26, 0, 23, 18, 0, 0, 0, 
		23, 35, 54, 0, 40, 39, 28, 51, 64, 44, 53, 58, 78, 67, 72, 
		96, 61, 37, 0, 95, 121, 98, 100, 103, 93, 101, 105, 108, 108, 115, 
		139, 93, 48, 41, 121, 97, 98, 95, 96, 100, 108, 113, 116, 120, 121, 
		145, 125, 82, 82, 96, 98, 103, 99, 98, 106, 120, 125, 129, 130, 143, 
		141, 127, 122, 92, 101, 102, 102, 98, 94, 105, 116, 111, 100, 129, 142, 
		
		0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 6, 4, 0, 0, 
		0, 0, 0, 0, 0, 15, 1, 4, 0, 19, 13, 13, 13, 4, 0, 
		0, 6, 0, 0, 0, 15, 0, 10, 13, 37, 20, 21, 0, 9, 5, 
		0, 24, 0, 0, 0, 19, 18, 8, 5, 43, 10, 13, 1, 0, 20, 
		20, 41, 0, 44, 56, 43, 27, 9, 1, 42, 35, 6, 15, 0, 8, 
		28, 44, 0, 0, 59, 41, 24, 21, 0, 68, 21, 7, 23, 11, 5, 
		37, 21, 17, 0, 37, 43, 42, 20, 8, 64, 18, 9, 15, 22, 5, 
		41, 48, 24, 13, 24, 65, 17, 19, 7, 38, 12, 7, 25, 16, 2, 
		43, 61, 3, 38, 8, 28, 17, 12, 33, 4, 22, 0, 10, 8, 0, 
		44, 51, 10, 53, 29, 21, 46, 32, 20, 14, 0, 11, 25, 16, 3, 
		64, 53, 15, 94, 26, 38, 52, 49, 20, 14, 24, 26, 29, 31, 19, 
		64, 61, 47, 80, 17, 18, 32, 32, 22, 24, 26, 30, 33, 32, 31, 
		20, 52, 74, 46, 18, 30, 27, 26, 23, 26, 33, 37, 34, 36, 47, 
		26, 30, 78, 24, 16, 34, 24, 28, 30, 33, 29, 31, 28, 44, 22, 
		24, 32, 22, 39, 14, 25, 26, 28, 32, 34, 26, 31, 50, 37, 16, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 12, 0, 0, 0, 18, 12, 12, 11, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 14, 12, 14, 0, 0, 0, 4, 0, 
		0, 42, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
		0, 3, 0, 20, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 19, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 6, 
		0, 0, 0, 0, 15, 5, 0, 0, 0, 26, 0, 0, 6, 0, 0, 
		0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 4, 0, 0, 
		0, 0, 0, 27, 0, 0, 19, 0, 0, 0, 0, 9, 15, 5, 0, 
		0, 0, 0, 31, 0, 0, 0, 0, 0, 9, 23, 15, 14, 5, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 14, 0, 3, 0, 0, 0, 0, 0, 0, 
		0, 3, 0, 0, 0, 0, 0, 17, 17, 0, 0, 9, 0, 11, 0, 
		0, 0, 0, 0, 0, 17, 0, 26, 0, 0, 0, 0, 0, 0, 0, 
		48, 0, 26, 58, 0, 50, 0, 1, 0, 35, 0, 16, 0, 0, 22, 
		118, 0, 38, 22, 0, 69, 0, 4, 0, 0, 21, 39, 0, 5, 15, 
		144, 0, 23, 0, 0, 0, 0, 19, 0, 0, 23, 8, 0, 0, 6, 
		92, 0, 78, 0, 24, 0, 47, 0, 0, 0, 0, 0, 0, 0, 23, 
		39, 0, 63, 0, 34, 31, 0, 0, 8, 0, 0, 26, 0, 0, 0, 
		0, 0, 0, 0, 0, 77, 34, 0, 34, 0, 15, 10, 0, 0, 1, 
		0, 4, 0, 0, 0, 14, 0, 0, 30, 19, 0, 0, 0, 0, 0, 
		0, 0, 43, 0, 0, 47, 0, 0, 3, 3, 0, 0, 0, 0, 2, 
		9, 0, 60, 0, 89, 0, 0, 0, 1, 0, 0, 0, 0, 11, 1, 
		9, 0, 30, 0, 27, 6, 3, 0, 2, 0, 3, 0, 7, 0, 0, 
		12, 0, 1, 0, 10, 0, 1, 9, 0, 0, 1, 12, 0, 0, 13, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 78, 0, 0, 0, 16, 27, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 3, 4, 0, 8, 
		0, 52, 0, 0, 9, 7, 24, 0, 8, 0, 0, 0, 0, 0, 0, 
		2, 50, 0, 0, 92, 33, 0, 0, 0, 23, 0, 0, 10, 10, 0, 
		0, 7, 0, 0, 0, 0, 31, 0, 12, 68, 0, 0, 0, 4, 19, 
		0, 3, 0, 0, 0, 42, 0, 14, 0, 41, 0, 0, 0, 12, 0, 
		0, 2, 0, 8, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
		0, 0, 0, 24, 0, 0, 0, 12, 1, 0, 0, 0, 0, 6, 12, 
		0, 0, 0, 21, 0, 0, 14, 37, 0, 0, 0, 0, 26, 21, 0, 
		18, 0, 0, 62, 115, 23, 32, 0, 0, 10, 14, 50, 24, 0, 0, 
		0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
		0, 0, 6, 0, 0, 0, 0, 0, 0, 1, 7, 6, 0, 0, 18, 
		0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 9, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 15, 13, 0, 0, 31, 4, 0, 
		
		46, 49, 50, 48, 46, 42, 53, 59, 47, 26, 18, 26, 35, 41, 44, 
		45, 53, 50, 49, 48, 25, 30, 30, 19, 0, 0, 0, 0, 23, 36, 
		11, 29, 52, 54, 53, 24, 20, 0, 0, 0, 0, 0, 0, 0, 26, 
		0, 0, 41, 46, 31, 12, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
		0, 0, 26, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 30, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 7, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 26, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 17, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 11, 0, 10, 0, 25, 10, 0, 0, 0, 
		10, 0, 0, 0, 0, 0, 37, 14, 0, 0, 46, 35, 51, 0, 0, 
		115, 0, 0, 0, 8, 0, 39, 28, 20, 0, 72, 13, 50, 22, 0, 
		115, 0, 28, 0, 55, 10, 71, 52, 36, 0, 43, 68, 19, 58, 0, 
		55, 8, 41, 0, 0, 16, 87, 59, 88, 0, 78, 74, 1, 43, 27, 
		49, 75, 0, 69, 0, 0, 63, 58, 99, 0, 99, 57, 3, 6, 37, 
		42, 91, 11, 50, 0, 0, 94, 27, 57, 0, 65, 68, 0, 5, 12, 
		73, 33, 97, 0, 11, 0, 40, 36, 0, 31, 0, 65, 0, 0, 0, 
		46, 27, 142, 0, 71, 0, 0, 79, 0, 26, 66, 16, 0, 0, 2, 
		0, 28, 129, 0, 157, 58, 0, 64, 92, 54, 19, 15, 3, 4, 31, 
		0, 1, 65, 0, 159, 78, 23, 29, 46, 34, 35, 31, 37, 34, 48, 
		56, 0, 0, 71, 149, 40, 44, 36, 39, 34, 33, 35, 42, 41, 36, 
		74, 33, 0, 161, 69, 30, 54, 39, 32, 34, 37, 43, 52, 22, 64, 
		82, 44, 18, 59, 44, 17, 33, 42, 33, 45, 56, 34, 11, 80, 102, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		3, 0, 2, 0, 4, 36, 10, 0, 0, 0, 18, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 1, 10, 9, 0, 0, 
		4, 23, 0, 0, 0, 0, 21, 14, 0, 0, 0, 0, 0, 0, 0, 
		45, 49, 11, 42, 79, 57, 0, 0, 0, 24, 21, 18, 1, 14, 0, 
		0, 0, 7, 0, 0, 0, 14, 15, 0, 46, 0, 0, 0, 7, 29, 
		30, 0, 0, 0, 0, 23, 0, 5, 0, 1, 0, 0, 0, 16, 12, 
		26, 0, 36, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		11, 0, 0, 8, 1, 0, 0, 0, 17, 0, 0, 0, 0, 8, 27, 
		0, 0, 0, 9, 0, 0, 12, 34, 0, 0, 0, 0, 21, 13, 0, 
		0, 0, 0, 58, 123, 85, 10, 0, 0, 0, 20, 46, 13, 0, 0, 
		0, 0, 29, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 5, 0, 0, 0, 0, 0, 0, 2, 7, 9, 0, 0, 15, 
		0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 5, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 14, 10, 0, 0, 38, 9, 0, 
		
		3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 15, 6, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 2, 34, 0, 0, 0, 8, 0, 0, 
		31, 15, 0, 0, 0, 68, 9, 11, 0, 0, 0, 0, 0, 17, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 21, 0, 0, 1, 
		0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 22, 
		29, 0, 0, 55, 53, 25, 0, 0, 0, 0, 21, 13, 0, 0, 0, 
		0, 5, 8, 0, 21, 0, 11, 0, 0, 0, 8, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 13, 60, 40, 0, 17, 3, 5, 0, 20, 0, 
		0, 0, 6, 0, 0, 60, 0, 0, 0, 12, 34, 50, 18, 0, 0, 
		5, 5, 0, 0, 3, 18, 0, 0, 20, 47, 40, 0, 0, 0, 0, 
		0, 0, 5, 0, 0, 0, 4, 41, 6, 0, 0, 0, 0, 0, 0, 
		79, 13, 0, 0, 111, 58, 43, 39, 6, 0, 0, 0, 0, 0, 0, 
		0, 63, 0, 42, 62, 0, 1, 0, 0, 0, 0, 0, 5, 3, 0, 
		0, 0, 64, 54, 3, 0, 0, 0, 0, 0, 5, 14, 0, 0, 56, 
		3, 0, 12, 50, 22, 23, 23, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		others=>0 );
END gold_package;
